/** 
 * 增加闹钟功能，最长闹铃时间为1分钟。闹钟的闹铃时刻可任意设置（只要求对时、分设置）。
 * 设置一个停止闹铃的按键，可以停止闹铃输出。 
 */

 module alarm