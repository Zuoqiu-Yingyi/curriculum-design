/* 菜单 */
module menu(
   input [1:0] FUN,
   
)